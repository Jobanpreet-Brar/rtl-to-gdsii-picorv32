

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO asic_top 
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 2.6968 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1124 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.0652 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 27.9676 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 105.45 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.13346 LAYER Via45 ;
  END clk
  PIN resetn 
    ANTENNAPARTIALMETALAREA 27.6168 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 104.749 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4914 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 106.067 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 405.879 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.2704 LAYER Via34 ;
    ANTENNAMAXCUTCAR 3.05397 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 23.9828 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 90.0576 LAYER Metal4 ;
    ANTENNAGATEAREA 3.6522 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 112.634 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 430.537 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAMAXCUTCAR 4.00841 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 32.5516 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 123.628 LAYER Metal5 ;
    ANTENNAGATEAREA 9.9486 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 115.906 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 442.964 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 5.05421 LAYER Via56 ;
  END resetn
  PIN mem_valid 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 6.4568 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.7404 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5112 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 226.016 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 858.528 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 2.60802 LAYER Via34 ;
  END mem_valid
  PIN mem_instr 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 7.7352 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.3832 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 33.8192 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 131.028 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.804762 LAYER Via34 ;
  END mem_instr
  PIN mem_ready 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 0.623 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3108 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 36.0352 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 162.301 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6156 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 83.5023 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 359.8 LAYER Metal6 ;
  END mem_ready
  PIN mem_addr[31] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 129.205 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 489.381 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal6 ; 
    ANTENNAPARTIALMETALAREA 25.506 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 114.919 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 126.683 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 555.34 LAYER Metal6 ;
  END mem_addr[31]
  PIN mem_addr[30] 
    ANTENNAPARTIALMETALAREA 3.0368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2996 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 1.3496 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.406 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 128.079 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 484.971 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 536.216 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 2034.15 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[30]
  PIN mem_addr[29] 
    ANTENNAPARTIALMETALAREA 11.5696 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 43.7992 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 4.3808 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.6844 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 116.93 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 442.762 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 487.045 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1846.04 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[29]
  PIN mem_addr[28] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 131.114 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 496.758 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 593.772 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 2252.04 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[28]
  PIN mem_addr[27] 
    ANTENNAPARTIALMETALAREA 5.6616 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.73 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 10.8504 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 40.9796 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 122.571 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 463.973 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal6 ; 
    ANTENNAPARTIALMETALAREA 33.0107 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 148.639 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 161.239 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 708.16 LAYER Metal6 ;
  END mem_addr[27]
  PIN mem_addr[26] 
    ANTENNAPARTIALMETALAREA 6.3112 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.8924 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 11.5938 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 43.7674 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 122.275 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 462.997 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 605.016 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 2293.43 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[26]
  PIN mem_addr[25] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.304 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 132.199 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 501.062 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 594.365 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 2255.07 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[25]
  PIN mem_addr[24] 
    ANTENNAPARTIALMETALAREA 3.948 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.946 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 14.0844 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 53.2226 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 63.5502 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 240.535 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal6 ; 
    ANTENNAPARTIALMETALAREA 12.6932 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 57.2616 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 385.68 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 1498.26 LAYER Metal6 ;
  END mem_addr[24]
  PIN mem_addr[23] 
    ANTENNAPARTIALMETALAREA 5.7528 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.5816 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 3.3012 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7942 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 125.785 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 476.088 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 542.263 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 2056.99 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[23]
  PIN mem_addr[22] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.2912 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3992 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 0.609 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2578 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal6 ; 
    ANTENNAPARTIALMETALAREA 3.8228 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 17.3448 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 570.53 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 2173.69 LAYER Metal6 ;
  END mem_addr[22]
  PIN mem_addr[21] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 125.195 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 474.202 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal6 ; 
    ANTENNAPARTIALMETALAREA 29.6376 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 133.511 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 144.591 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 634.377 LAYER Metal6 ;
  END mem_addr[21]
  PIN mem_addr[20] 
    ANTENNAPARTIALMETALAREA 3.024 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.448 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 4.4496 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.748 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 127.994 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 484.844 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 546.622 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 2071.58 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 2.14603 LAYER Via56 ;
  END mem_addr[20]
  PIN mem_addr[19] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 115.825 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 438.681 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 581.227 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 2204.55 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[19]
  PIN mem_addr[18] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 16.6026 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 62.805 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal6 ; 
    ANTENNAPARTIALMETALAREA 8.9972 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 40.6296 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 519.08 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 1993.22 LAYER Metal6 ;
  END mem_addr[18]
  PIN mem_addr[17] 
    ANTENNAPARTIALMETALAREA 4.844 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.338 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 5.0768 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.1224 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 86.156 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 326.459 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 386.194 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1465.03 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 2.14603 LAYER Via56 ;
  END mem_addr[17]
  PIN mem_addr[16] 
    ANTENNAPARTIALMETALAREA 2.9848 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2996 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.304 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 85.2504 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 323.13 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 403.527 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1531.83 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[16]
  PIN mem_addr[15] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.304 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 97.3616 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 368.88 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 402.572 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1527.03 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[15]
  PIN mem_addr[14] 
    ANTENNAPARTIALMETALAREA 6.5072 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.6344 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 4.164 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6668 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 83.4848 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 316.346 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 366.673 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1393.35 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 2.14603 LAYER Via56 ;
  END mem_addr[14]
  PIN mem_addr[13] 
    ANTENNAPARTIALMETALAREA 4.7936 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.444 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 2.6292 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.2502 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 79.9136 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 302.63 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 336.111 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1275.83 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[13]
  PIN mem_addr[12] 
    ANTENNAPARTIALMETALAREA 5.5832 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1364 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 2.0176 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.738 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 73.5148 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 278.398 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 325.835 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1236.5 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[12]
  PIN mem_addr[11] 
    ANTENNAPARTIALMETALAREA 6.1376 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.2352 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 1.5992 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9572 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 75.6336 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 286.624 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 319.349 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1211.98 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 2.14603 LAYER Via56 ;
  END mem_addr[11]
  PIN mem_addr[10] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 78.2096 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 296.376 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 331.365 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1258.25 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[10]
  PIN mem_addr[9] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.9452 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6782 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 59.7688 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 226.564 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 291.099 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1105.81 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[9]
  PIN mem_addr[8] 
    ANTENNAPARTIALMETALAREA 0.6344 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2048 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.8904 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6676 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 13.4248 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 50.9224 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 93.7938 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 358.087 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_addr[8]
  PIN mem_addr[7] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 16.6432 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.0064 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 89.8542 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 340.84 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.07302 LAYER Via34 ;
  END mem_addr[7]
  PIN mem_addr[6] 
    ANTENNAPARTIALMETALAREA 4.1048 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.5396 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.0696 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.738 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 69.1653 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 265.084 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 1.60952 LAYER Via45 ;
  END mem_addr[6]
  PIN mem_addr[5] 
    ANTENNAPARTIALMETALAREA 4.5284 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9388 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 13.9344 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 52.8516 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 98.8764 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 378.109 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 1.34127 LAYER Via45 ;
  END mem_addr[5]
  PIN mem_addr[4] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 8.5136 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.6268 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 38.2081 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 149.241 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.804762 LAYER Via34 ;
  END mem_addr[4]
  PIN mem_addr[3] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 8.8592 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.8352 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 49.7637 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 195.595 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.07302 LAYER Via34 ;
  END mem_addr[3]
  PIN mem_addr[2] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 10.8768 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 41.2764 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 51.647 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 199.465 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.07302 LAYER Via34 ;
  END mem_addr[2]
  PIN mem_wdata[31] 
    ANTENNAPARTIALMETALAREA 0.6344 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2048 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 4.1848 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9424 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3993 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 62.1069 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 237.312 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.18507 LAYER Via56 ;
  END mem_wdata[31]
  PIN mem_wdata[30] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 5.4548 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5004 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 8.1984 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 31.3336 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3993 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 67.1362 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 256.465 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.18507 LAYER Via56 ;
  END mem_wdata[30]
  PIN mem_wdata[29] 
    ANTENNAPARTIALMETALAREA 8.26 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.27 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 17.6812 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 66.5892 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3993 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 51.2534 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 195.462 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.846481 LAYER Via45 ;
  END mem_wdata[29]
  PIN mem_wdata[28] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 11.1776 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.612 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3993 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 30.9269 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 119.379 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.507889 LAYER Via34 ;
  END mem_wdata[28]
  PIN mem_wdata[27] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 3.569 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3878 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 10.64 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.5768 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3993 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 51.5214 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 197.731 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.18507 LAYER Via56 ;
  END mem_wdata[27]
  PIN mem_wdata[26] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 14 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 53 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3993 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 45.0466 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 171.596 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.507889 LAYER Via34 ;
  END mem_wdata[26]
  PIN mem_wdata[25] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 6.6544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.2916 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3993 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 21.0676 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 82.0551 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.507889 LAYER Via34 ;
  END mem_wdata[25]
  PIN mem_wdata[24] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.2912 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3992 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 3.4328 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.2924 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3993 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 34.6078 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 133.568 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.18507 LAYER Via56 ;
  END mem_wdata[24]
  PIN mem_wdata[23] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 15.3456 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 58.194 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.36 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 62.4331 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 238.971 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.50222 LAYER Via56 ;
  END mem_wdata[23]
  PIN mem_wdata[22] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 20.2832 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 76.7864 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.36 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 63.1164 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 240.178 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.751111 LAYER Via34 ;
  END mem_wdata[22]
  PIN mem_wdata[21] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 13.8712 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 52.5124 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.36 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 52.7119 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 203.019 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.751111 LAYER Via34 ;
  END mem_wdata[21]
  PIN mem_wdata[20] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 22.5008 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 85.1816 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.36 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 67.9401 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 258.243 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.751111 LAYER Via34 ;
  END mem_wdata[20]
  PIN mem_wdata[19] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 5.848 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.2388 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.36 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 55.3394 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 211.176 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.31444 LAYER Via56 ;
  END mem_wdata[19]
  PIN mem_wdata[18] 
    ANTENNAPARTIALMETALAREA 3.0368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.2996 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 4.224 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0908 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 10.8248 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 41.2764 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.36 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 59.1008 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 225.809 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.50222 LAYER Via56 ;
  END mem_wdata[18]
  PIN mem_wdata[17] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 22.5976 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 85.3512 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.36 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 65.9179 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 250.587 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.751111 LAYER Via34 ;
  END mem_wdata[17]
  PIN mem_wdata[16] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 16.88 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 64.0028 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.36 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 84.1328 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 320.179 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.50222 LAYER Via56 ;
  END mem_wdata[16]
  PIN mem_wdata[15] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 24.1589 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 93.6754 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.536508 LAYER Via34 ;
  END mem_wdata[15]
  PIN mem_wdata[14] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 5.6072 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.3272 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 99.8692 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 381.432 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 2.14603 LAYER Via56 ;
  END mem_wdata[14]
  PIN mem_wdata[13] 
    ANTENNAPARTIALMETALAREA 0.6344 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2048 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 2.3016 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.01 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 3.3896 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.932 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 89.4065 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 339.915 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 2.14603 LAYER Via56 ;
  END mem_wdata[13]
  PIN mem_wdata[12] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 6.4288 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.6344 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 36.8859 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 142.637 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.804762 LAYER Via34 ;
  END mem_wdata[12]
  PIN mem_wdata[11] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 8.7544 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.9448 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 49.5486 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 189.538 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.07302 LAYER Via34 ;
  END mem_wdata[11]
  PIN mem_wdata[10] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 7.5504 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.6836 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 35.5304 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 137.506 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.804762 LAYER Via34 ;
  END mem_wdata[10]
  PIN mem_wdata[9] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 38.52 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 165.394 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 0.804762 LAYER Via34 ;
  END mem_wdata[9]
  PIN mem_wdata[8] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 7.1936 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.136 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 46.8843 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 179.948 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.07302 LAYER Via34 ;
  END mem_wdata[8]
  PIN mem_wdata[7] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.6584 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.9496 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 39.1103 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 150.739 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.56481 LAYER Via34 ;
  END mem_wdata[7]
  PIN mem_wdata[6] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.5128 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3984 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 35.4807 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 136.998 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.56481 LAYER Via34 ;
  END mem_wdata[6]
  PIN mem_wdata[5] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.6848 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2464 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 36.4205 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 140.556 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 2.08642 LAYER Via34 ;
  END mem_wdata[5]
  PIN mem_wdata[4] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 2.9456 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.448 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 38.2909 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 146.118 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 2.08642 LAYER Via34 ;
  END mem_wdata[4]
  PIN mem_wdata[3] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 7.2088 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.3904 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 63.6119 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 241.976 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 2.08642 LAYER Via34 ;
  END mem_wdata[3]
  PIN mem_wdata[2] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.6456 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.098 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 34.1721 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 133.563 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.04321 LAYER Via34 ;
  END mem_wdata[2]
  PIN mem_wdata[1] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 4.7936 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.444 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 44.9761 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 172.945 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 2.08642 LAYER Via34 ;
  END mem_wdata[1]
  PIN mem_wdata[0] 
    ANTENNADIFFAREA 0.5176 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 3.276 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6988 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 39.6304 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 151.189 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 2.08642 LAYER Via34 ;
  END mem_wdata[0]
  PIN mem_wstrb[3] 
    ANTENNAPARTIALMETALAREA 3.8808 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.6916 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 22.6566 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 85.648 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3633 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 94.0149 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 358.206 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.930361 LAYER Via45 ;
  END mem_wstrb[3]
  PIN mem_wstrb[2] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 3.3896 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 12.932 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3633 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 97.6764 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 371.598 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.3025 LAYER Via56 ;
  END mem_wstrb[2]
  PIN mem_wstrb[1] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 1.4424 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3636 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 4.9518 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.6984 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal6 ; 
    ANTENNAPARTIALMETALAREA 35.2476 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 158.756 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3024 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 154.594 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 670.633 LAYER Metal6 ;
  END mem_wstrb[1]
  PIN mem_wstrb[0] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNADIFFAREA 0.5176 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 6.2176 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.638 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1368 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 244.887 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 931.336 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 3.95322 LAYER Via56 ;
  END mem_wstrb[0]
  PIN mem_rdata[31] 
    ANTENNAPARTIALMETALAREA 14.78 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.756 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 21.4456 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 81.6836 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5738 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 139.533 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 529.063 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 6.04448 LAYER Via56 ;
  END mem_rdata[31]
  PIN mem_rdata[30] 
    ANTENNAPARTIALMETALAREA 12.1984 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 46.2796 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 2.6104 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9852 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 74.9082 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 284.016 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAMAXCUTCAR 5.21605 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 12.8562 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 48.6222 LAYER Metal5 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 174.107 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 659.188 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 7.21605 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 52.7438 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 237.125 LAYER Metal6 ;
    ANTENNAGATEAREA 1.6524 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 206.027 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 802.691 LAYER Metal6 ;
  END mem_rdata[30]
  PIN mem_rdata[29] 
    ANTENNAPARTIALMETALAREA 8.3552 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.6304 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.5016 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.802 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 23.415 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 88.5948 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 67.102 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 255.33 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 4.70225 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 56.1344 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 252.747 LAYER Metal6 ;
    ANTENNAGATEAREA 1.6524 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 111.952 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 451.117 LAYER Metal6 ;
  END mem_rdata[29]
  PIN mem_rdata[28] 
    ANTENNAPARTIALMETALAREA 5.9808 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6416 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 7.244 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.3268 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 91.8436 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 348.38 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3899 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 140.295 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 534.511 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 4.17284 LAYER Via56 ;
  END mem_rdata[28]
  PIN mem_rdata[27] 
    ANTENNAPARTIALMETALAREA 8.1984 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.0368 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.5016 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.802 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 24.6318 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 93.0044 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 64.5963 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 249.012 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 3.65904 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 42.886 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 193.129 LAYER Metal6 ;
    ANTENNAGATEAREA 1.6524 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 92.979 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 373.401 LAYER Metal6 ;
  END mem_rdata[27]
  PIN mem_rdata[26] 
    ANTENNAPARTIALMETALAREA 7.472 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.09 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.6176 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.438 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 21.8414 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 82.9344 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 87.7658 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 333.177 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 5.74546 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 55.6795 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 250.648 LAYER Metal6 ;
    ANTENNAGATEAREA 1.6524 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 125.271 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 501.312 LAYER Metal6 ;
  END mem_rdata[26]
  PIN mem_rdata[25] 
    ANTENNAPARTIALMETALAREA 7.6008 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.5776 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 5.5862 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.2 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 77.1609 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 292.469 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 5.25454 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 50.146 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 225.799 LAYER Metal6 ;
    ANTENNAGATEAREA 1.3899 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 160.316 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 636.219 LAYER Metal6 ;
  END mem_rdata[25]
  PIN mem_rdata[24] 
    ANTENNAPARTIALMETALAREA 12.992 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.184 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 4.3352 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5148 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 80.0934 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 303.646 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAMAXCUTCAR 5.21605 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 10.4398 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 39.4744 LAYER Metal5 ;
    ANTENNAGATEAREA 0.4896 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 101.416 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 384.272 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 5.74546 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 29.6948 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 133.769 LAYER Metal6 ;
    ANTENNAGATEAREA 1.6131 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 119.825 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 467.198 LAYER Metal6 ;
  END mem_rdata[24]
  PIN mem_rdata[23] 
    ANTENNAPARTIALMETALAREA 5.1632 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8432 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 2.3424 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.9676 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 58.4672 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 221.54 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1598 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 136.984 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 518.854 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 4.17284 LAYER Via56 ;
  END mem_rdata[23]
  PIN mem_rdata[22] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.4228 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8974 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 4.7238 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 17.6384 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 15.782 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 71.1612 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.218 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 121 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 469.416 LAYER Metal6 ;
  END mem_rdata[22]
  PIN mem_rdata[21] 
    ANTENNAPARTIALMETALAREA 7.5392 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.6412 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.5548 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9504 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 31.4986 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 119.494 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3816 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 171.729 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 651.954 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 6.9385 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 8.5044 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 38.412 LAYER Metal6 ;
    ANTENNAGATEAREA 1.11 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 179.391 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 686.56 LAYER Metal6 ;
  END mem_rdata[21]
  PIN mem_rdata[20] 
    ANTENNAPARTIALMETALAREA 11.7264 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.3928 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 12.9116 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 48.9826 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 181.251 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 685.851 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAMAXCUTCAR 6.25926 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 23.9024 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 90.5876 LAYER Metal5 ;
    ANTENNAGATEAREA 1.2544 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 200.306 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 758.067 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 6.25926 LAYER Via56 ;
  END mem_rdata[20]
  PIN mem_rdata[19] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.6316 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.491 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 33.1702 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 125.822 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 129.613 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 493.117 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 4.70225 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 13.802 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 62.2512 LAYER Metal6 ;
    ANTENNAGATEAREA 1.2502 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 140.653 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 542.91 LAYER Metal6 ;
  END mem_rdata[19]
  PIN mem_rdata[18] 
    ANTENNAPARTIALMETALAREA 13.1264 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.9896 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.304 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 17.0928 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 65.1052 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2544 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 83.2906 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 317.924 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 6.25926 LAYER Via56 ;
  END mem_rdata[18]
  PIN mem_rdata[17] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 1.7178 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.4554 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 15.8964 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 71.676 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2502 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 89.829 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 350.206 LAYER Metal6 ;
  END mem_rdata[17]
  PIN mem_rdata[16] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 1.232 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9608 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 2.8394 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5046 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 18.4924 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 83.358 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2544 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 76.7383 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 303.058 LAYER Metal6 ;
  END mem_rdata[16]
  PIN mem_rdata[15] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 1.218 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.9078 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 34.3144 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 130.104 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.489 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 54.9169 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 209.14 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.29929 LAYER Via56 ;
  END mem_rdata[15]
  PIN mem_rdata[14] 
    ANTENNAPARTIALMETALAREA 0.6344 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2048 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 37.4238 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 141.531 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7606 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 64.2698 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 244.281 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 1.80291 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 29.0824 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 131.155 LAYER Metal6 ;
    ANTENNAGATEAREA 1.4848 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 135.61 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 528.438 LAYER Metal6 ;
  END mem_rdata[14]
  PIN mem_rdata[13] 
    ANTENNAPARTIALMETALAREA 3.1936 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8932 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.7336 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.074 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 37.1786 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 140.503 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7606 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 57.4817 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 221.951 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 1.16073 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 19.0996 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 86.0904 LAYER Metal6 ;
    ANTENNAGATEAREA 1.4848 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 130.5 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 504.368 LAYER Metal6 ;
  END mem_rdata[13]
  PIN mem_rdata[12] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 1.0054 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5616 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 4.8084 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.78 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3902 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 120.208 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 459.646 LAYER Metal6 ;
  END mem_rdata[12]
  PIN mem_rdata[11] 
    ANTENNAPARTIALMETALAREA 3.1416 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8932 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 4.7112 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9352 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 19.2074 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 72.4616 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 27.0612 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 121.473 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4442 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 68.5953 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 273.733 LAYER Metal6 ;
  END mem_rdata[11]
  PIN mem_rdata[10] 
    ANTENNAPARTIALMETALAREA 29.3848 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 111.639 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.72 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 56.2722 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 215.725 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAMAXCUTCAR 1.31444 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 19.3668 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 73.0234 LAYER Metal4 ;
    ANTENNAGATEAREA 1.0842 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 74.1349 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 283.077 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAMAXCUTCAR 1.43914 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 59.6512 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 226.416 LAYER Metal5 ;
    ANTENNAGATEAREA 1.4442 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 115.439 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 439.853 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.50222 LAYER Via56 ;
  END mem_rdata[10]
  PIN mem_rdata[9] 
    ANTENNAPARTIALMETALAREA 11.6536 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.1172 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 1.756 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5508 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 68.484 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 259.954 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4848 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 69.7217 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 267.179 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.50222 LAYER Via56 ;
  END mem_rdata[9]
  PIN mem_rdata[8] 
    ANTENNAPARTIALMETALAREA 4.8328 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2956 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.8152 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9892 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 33.8534 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 128.112 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7606 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 50.5006 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 193.241 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAMAXCUTCAR 1.84301 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 19.2316 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 86.6844 LAYER Metal6 ;
    ANTENNAGATEAREA 1.489 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 141.525 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 547.12 LAYER Metal6 ;
  END mem_rdata[8]
  PIN mem_rdata[7] 
    ANTENNAPARTIALMETALAREA 0.6344 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.2048 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.5768 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4804 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 20.712 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 78.6096 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.063 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 56.9473 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 217.72 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.78836 LAYER Via56 ;
  END mem_rdata[7]
  PIN mem_rdata[6] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 0.1064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6996 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 1.3482 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.0562 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.2592 LAYER Via56 ;
    ANTENNAPARTIALMETALAREA 9.3756 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 42.3324 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.063 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 64.6163 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 251.819 LAYER Metal6 ;
  END mem_rdata[6]
  PIN mem_rdata[5] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 5.82 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1328 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 22.9096 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 87.026 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0224 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 45.5391 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 174.422 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.47351 LAYER Via56 ;
  END mem_rdata[5]
  PIN mem_rdata[4] 
    ANTENNAPARTIALMETALAREA 0.252 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.954 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 2.4724 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.6566 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 28.4664 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 107.866 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1206 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 57.2718 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 218.049 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 0.804633 LAYER Via56 ;
  END mem_rdata[4]
  PIN mem_rdata[3] 
    ANTENNAPARTIALMETALAREA 5.0568 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.1436 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 8.9688 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.8564 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 23.7608 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 90.2484 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1206 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 34.2746 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 131.527 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.50222 LAYER Via56 ;
  END mem_rdata[3]
  PIN mem_rdata[2] 
    ANTENNAPARTIALMETALAREA 0.4368 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6536 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0676 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 5.2948 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.3414 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via45 ;
    ANTENNAPARTIALMETALAREA 30.7304 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 116.536 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1206 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 42.5179 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 162.147 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.87778 LAYER Via56 ;
  END mem_rdata[2]
  PIN mem_rdata[1] 
    ANTENNAPARTIALMETALAREA 26.0976 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 99.1948 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8955 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 39.5303 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 155.053 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAMAXCUTCAR 2.12759 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 3.4808 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0804 LAYER Metal4 ;
    ANTENNAGATEAREA 1.2555 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 42.3027 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 165.472 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 2.12759 LAYER Via45 ;
  END mem_rdata[1]
  PIN mem_rdata[0] 
    ANTENNAPARTIALMETALAREA 11.8288 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 44.8804 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER Via34 ;
    ANTENNAPARTIALMETALAREA 8.8584 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.5384 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2961 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 51.4446 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 196.185 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 3.10925 LAYER Via45 ;
  END mem_rdata[0]
  PIN trap 
    ANTENNADIFFAREA 0.72 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 16.1408 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 61.2044 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 96.8265 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 367.859 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.25185 LAYER Via34 ;
  END trap
END asic_top

END LIBRARY
